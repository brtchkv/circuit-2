`timescale 1ns / 1ps

module mult(
    input clk,
    input rst,
    input start,
    input [7:0] a,
    input [7:0] b,
    output wire ready,
    output wire busy,
    output reg [15:0] y
);

localparam IDLE =      1'b0;
localparam WORK =      1'b1;

reg [2:0] ctr;
wire [2:0] end_step;
wire [7:0] part_sum;
wire [15:0] shifted_part_sum;
reg [15:0] part_res;

reg state;
reg ready_in;

assign part_sum = a & { 8{ b[ctr] }};
assign shifted_part_sum = part_sum << ctr;
assign end_step = (ctr == 3'h7);
assign busy = state;
assign ready = ready_in;

always @(posedge clk)
    if (rst) begin
        ctr <= 0;
        part_res <= 0;
        y <= 0;
        state <= IDLE;
        ready_in <= 1;
    end else begin
        case (state)
            IDLE: 
                if (ready && start) begin
                    state <= WORK;
                    ctr <= 0;
                    part_res <= 0;
                    ready_in <= 0;
                end
            WORK:
                begin
                    if (end_step) begin
                        state <= IDLE;
                        y <= part_res;
                    end
                    
                    part_res <= part_res + shifted_part_sum;
                    ctr <= ctr + 1;
                end
        endcase
    end
endmodule